module LALU()

endmodule;