module VGA ();

endmodule