module VGA (
    input CLOCK_50,

    input charWr,
    input [23:0] charWrFgColor,
    input [23:0] charWrBgColor,
    input [7:0] charWrCode,
    input [5:0] charWrX,
    input [4:0] charWrY,

    output [7:0] VGA_R, VGA_G, VGA_B,
    output VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, VGA_HS, VGA_VS
);
    integer i;
    /*********************
     **      CHARS      **
     *********************/
    reg [0:199] characters[0:255];

    initial
    begin
        for (i = 0; i < 256; i = i + 1) characters[0] = 200'b0;

    	characters[65] = 200'b00001100000001001000000100100000010010000001001000001000010000100001000011111100001000010001000000100100000010010000001001000000100100000010010000001001000000100000000000000000000000000000000000000000;
    	characters[66] = 200'b01111110000100000100010000001001000000100100000010010000001001000001000111111000010000010001000000100100000010010000001001000000100100000010010000010001111110000000000000000000000000000000000000000000;
    	characters[67] = 200'b00011111100010000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000001000000000011111100000000000000000000000000000000000000000;
    	characters[68] = 200'b01111110000100000100010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000010001111110000000000000000000000000000000000000000000;
    	characters[69] = 200'b00111111100100000000010000000001000000000100000000010000000001000000000111111110010000000001000000000100000000010000000001000000000100000000010000000000111111100000000000000000000000000000000000000000;
    	characters[70] = 200'b00111111100100000000010000000001000000000100000000010000000001111111100100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000000000000000000000000000000000000000000;
    	characters[71] = 200'b00011111100010000000010000000001000000000100000000010000000001000000000100000000010000111001000000100100000010010000001001000000100100000010001000001000011111100000000000000000000000000000000000000000;
    	characters[72] = 200'b01000000100100000010010000001001000000100100000010010000001001000000100111111110010000001001000000100100000010010000001001000000100100000010010000001001000000100000000000000000000000000000000000000000;
    	characters[73] = 200'b01111111100000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000001111111100000000000000000000000000000000000000000;
    	characters[74] = 200'b00011111100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100100000010010000010000111110000000000000000000000000000000000000000000;
    	characters[75] = 200'b01000000100100000010010000001001000001000100001000010000100001001100000111000000010010000001001100000100001000010000100001000001000100000010010000001001000000100000000000000000000000000000000000000000;
    	characters[76] = 200'b01000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001111111100000000000000000000000000000000000000000;
    	characters[77] = 200'b01100001100101001010010100101001001100100100110010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100000000000000000000000000000000000000000;
    	characters[78] = 200'b01100000100101000010010100001001010000100100100010010010001001001000100100010010010001001001000100100100010010010000101001000010100100001010010000101001000001100000000000000000000000000000000000000000;
    	characters[79] = 200'b00111111000100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001000111111000000000000000000000000000000000000000000;
    	characters[80] = 200'b01111110000100000100010000001001000000100100000010010000001001000001000111111000010000000001000000000100000000010000000001000000000100000000010000000001000000000000000000000000000000000000000000000000;
    	characters[81] = 200'b00011110000010000100010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010010001001000100100100001010001000010000011110100000000000000000000000000000000000000000;
    	characters[82] = 200'b01111110000100000100010000001001000000100100000010010000001001000001000111111000011000000001011000000100010000010000100001000001000100000100010000001001000000100000000000000000000000000000000000000000;
    	characters[83] = 200'b00011110000010000100010000001001000000100100000000010000000000100000000001111000000000010000000000100000000010000000001001000000100100000010001000010000011110000000000000000000000000000000000000000000;
    	characters[84] = 200'b01111111100000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000000000000000000000000000000000000000;
    	characters[85] = 200'b01000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010001000010000011110000000000000000000000000000000000000000000;
    	characters[86] = 200'b01000000100100000010010000001001000000100100000010010000001000100001000010000100001000010000100001000010000100000100100000010010000001001000000100100000001100000000000000000000000000000000000000000000;
    	characters[87] = 200'b01000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100110010010011001001010010100101001010010100101001100001100000000000000000000000000000000000000000;
    	characters[88] = 200'b01000000100100000010001000010000100001000001001000000100100000010010000000110000000011000000010010000001001000000100100000100001000010000100010000001001000000100000000000000000000000000000000000000000;
    	characters[89] = 200'b01000000100100000010001000010000100001000001001000000100100000010010000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000000000000000000000000000000000000000;
    	characters[90] = 200'b01111111100000000010000000010000000010000000001000000001000000000100000000100000000010000000010000000001000000001000000000100000000100000000010000000001111111100000000000000000000000000000000000000000;
    end

    reg vga_clk;                    // VGA runs at 25MHz
    always @(posedge CLOCK_50) begin
        vga_clk <= ~vga_clk;
    end

    /*********************
     **     COUNTER     **
     *********************/
    reg [9:0] hCount = 0;
    reg [9:0] vCount = 0;

    wire hDisp = hCount < 640;
    wire vDisp = vCount < 480;

    reg [5:0] charX = 0;
    reg [4:0] charY = 0;
    reg [3:0] charU = 0;
    reg [4:0] charV = 0;

    always @(posedge vga_clk)
    begin
    	// NEW LINE
    	if (hCount == 799)
    	begin
    		hCount <= 0;
    		charX <= 0;
    		charU <= 0;

    		// NEW FRAME
    		if (vCount == 524)
    		begin
    			vCount <= 0;
    			charY <= 0;
    			charV <= 0;
    		end
    		// MID FRAME
    		else
    		begin
    			vCount <= vCount + 1;

    			// END CHAR
    			if (charV == 19)
    			begin
    				charV <= 0;
    				charY <= charY + 1;
    			end
    			// MID CHAR
    			else
    			begin
    				charV <= charV + 1;
    			end
    		end
    	end
    	// MID LINE
    	else
    	begin
    		hCount <= hCount + 1;

    		// END CHAR
    		if (charU == 9)
    		begin
    			charU <= 0;
    			charX <= charX + 1;
    		end
    		// MID CHAR
    		else
    		begin
    			charU <= charU + 1;
    		end
    	end
    end


    wire [55:0] vramOut;
    RAM #(11, 56, "MLAB") vram (
        .clk(CLOCK_50),

        .address_a(charWrX + charWrY * 64),
        .wren_a(charWr),
        .data_a({charWrFgColor, charWrBgColor, charWrCode}),
        .rden_a(1'b0),
        .q_a(),

        .address_b(charX + charY * 64),
        .wren_b(1'b0),
        .data_b(32'b0),
        .rden_b(1'b1),
        .q_b(vramOut)
    );

    wire [199:0] character = characters[vramOut[7:0]];
    wire [23:0] color = character[charU + charV*10] ? vramOut[31:8] : vramOut[55:32];

    assign VGA_CLK = vga_clk;
    assign VGA_HS = ~(656 <= hCount && hCount < 752);
    assign VGA_VS = ~(490 <= vCount && vCount < 492);
    assign VGA_R = color[23:16];
    assign VGA_B = color[15:8];
    assign VGA_G = color[7:0];
    assign VGA_BLANK_N = ~(~hDisp || ~vDisp);
    assign VGA_SYNC_N = 1'b1;

endmodule