module VGA (
    input CLOCK_50,

    input charWr,
    input [23:0] charWrFgColor,
    input [23:0] charWrBgColor,
    input [7:0] charWrCode,
    input [7:0] charWrFlags,
    input [5:0] charWrX,
    input [4:0] charWrY,

    output [7:0] VGA_R, VGA_G, VGA_B,
    output VGA_CLK, VGA_SYNC_N, VGA_BLANK_N, VGA_HS, VGA_VS
);
    parameter H_VISIBLE = 640;
    parameter H_FPORCH = 16;
    parameter H_SYNC = 96;
    parameter H_BPORCH = 48;
    parameter H_BP_END = H_BPORCH - 1;
    parameter H_END = H_VISIBLE + H_FPORCH + H_SYNC + H_BPORCH - 1;

    parameter V_VISIBLE = 480;
    parameter V_FPORCH = 10;
    parameter V_SYNC = 2;
    parameter V_BPORCH = 33;
    parameter V_BP_END = V_BPORCH - 1;
    parameter V_END = V_VISIBLE + V_FPORCH + V_SYNC + V_BPORCH - 1;

	clock25 gen(.CLOCK_50(CLOCK_50), .CLOCK_25(VGA_CLK));

    integer i;
    /*********************
     **      CHARS      **
     *********************/
    reg [0:159] characters[0:255];
    reg [0:159] boldCharacters[0:255];
    reg [0:159] italicCharacters[0:255];
    reg [0:159] boldItalicCharacters[0:255];

    initial
    begin
        for (i = 0; i < 256; i = i + 1) begin
            characters[i] = 160'b0;
            boldCharacters[i] = 160'b0;
            italicCharacters[i] = 160'b0;
            boldItalicCharacters[i] = 160'b0;
        end

    	characters[65] = 160'b0000110000000100100000010010000001001000000100100000100001000010000100001111110000100001000100000010010000001001000000100100000010010000001001000000100100000010;
    	characters[66] = 160'b0111111000010000010001000000100100000010010000001001000000100100000100011111100001000001000100000010010000001001000000100100000010010000001001000001000111111000;
    	characters[67] = 160'b0001111110001000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000000100000000001111110;
    	characters[68] = 160'b0111111000010000010001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000001000111111000;
    	characters[69] = 160'b0011111110010000000001000000000100000000010000000001000000000100000000011111111001000000000100000000010000000001000000000100000000010000000001000000000011111110;
    	characters[70] = 160'b0011111110010000000001000000000100000000010000000001000000000111111110010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000;
    	characters[71] = 160'b0001111110001000000001000000000100000000010000000001000000000100000000010000000001000011100100000010010000001001000000100100000010010000001000100000100001111110;
    	characters[72] = 160'b0100000010010000001001000000100100000010010000001001000000100100000010011111111001000000100100000010010000001001000000100100000010010000001001000000100100000010;
    	characters[73] = 160'b0111111110000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000111111110;
    	characters[74] = 160'b0001111110000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010010000001001000001000011111000;
    	characters[75] = 160'b0100000010010000001001000000100100000100010000100001000010000100110000011100000001001000000100110000010000100001000010000100000100010000001001000000100100000010;
    	characters[76] = 160'b0100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000100000000010000000001000000000111111110;
    	characters[77] = 160'b0110000110010100101001010010100100110010010011001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010;
    	characters[78] = 160'b0110000010010100001001010000100101000010010010001001001000100100100010010001001001000100100100010010010001001001000010100100001010010000101001000010100100000110;
    	characters[79] = 160'b0011111100010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100011111100;
    	characters[80] = 160'b0111111000010000010001000000100100000010010000001001000000100100000100011111100001000000000100000000010000000001000000000100000000010000000001000000000100000000;
    	characters[81] = 160'b0001111000001000010001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001001000100100010010010000101000100001000001111010;
    	characters[82] = 160'b0111111000010000010001000000100100000010010000001001000000100100000100011111100001100000000101100000010001000001000010000100000100010000010001000000100100000010;
    	characters[83] = 160'b0001111000001000010001000000100100000010010000000001000000000010000000000111100000000001000000000010000000001000000000100100000010010000001000100001000001111000;
    	characters[84] = 160'b0111111110000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000;
    	characters[85] = 160'b0100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010000001000100001000001111000;
    	characters[86] = 160'b0100000010010000001001000000100100000010010000001001000000100010000100001000010000100001000010000100001000010000010010000001001000000100100000010010000000110000;
    	characters[87] = 160'b0100000010010000001001000000100100000010010000001001000000100100000010010000001001000000100100000010010011001001001100100101001010010100101001010010100110000110;
    	characters[88] = 160'b0100000010010000001000100001000010000100000100100000010010000001001000000011000000001100000001001000000100100000010010000010000100001000010001000000100100000010;
    	characters[89] = 160'b0100000010010000001000100001000010000100000100100000010010000001001000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000;
    	characters[90] = 160'b0111111110000000001000000001000000001000000000100000000100000000010000000010000000001000000001000000000100000000100000000010000000010000000001000000000111111110;

        boldCharacters[65] = 200'b0000110000000111100000110011000011001100001100110000110011000011111100011111111001100001100110000110011000011001100001100110000110011000011001100001100110000110;
        boldCharacters[66] = 200'b0111111000011111110001100001100110000110011000011001100001100111111110011111110001111111100110000110011000011001100001100110000110011000011001111111000111111000;
        boldCharacters[67] = 200'b0001111110001111111001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000000111111100001111110;
        boldCharacters[68] = 200'b0111111000011111110001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011001111111000111111000;
        boldCharacters[69] = 200'b0011111110011111111001100000000110000000011000000001100000000110000000011111111001111111100110000000011000000001100000000110000000011000000001111111100011111110;
        boldCharacters[70] = 200'b0011111110011111111001100000000110000000011000000001100000000111111110011111111001100000000110000000011000000001100000000110000000011000000001100000000110000000;
        boldCharacters[71] = 200'b0001111110001111111001100000000110000000011000000001100000000110000000011000000001100011100110001110011000011001100001100110000110011000011000111111100001111110;
        boldCharacters[72] = 200'b0110000110011000011001100001100110000110011000011001100001100110000110011111111001111111100110000110011000011001100001100110000110011000011001100001100110000110;
        boldCharacters[73] = 200'b0111111110011111111000011110000001111000000111100000011110000001111000000111100000011110000001111000000111100000011110000001111000000111100001111111100111111110;
        boldCharacters[74] = 200'b0001111110000111111000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110011000011001111111000011111000;
        boldCharacters[75] = 200'b0110000110011000011001100001100110001100011000110001101110000111110000011100000001111000000111110000011011100001100110000110001100011000011001100001100110000110;
        boldCharacters[76] = 200'b0110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000000011000000001111111100111111110;
        boldCharacters[77] = 200'b0110000110011100111001110011100111111110011111111001101101100110000110011000011001100001100110000110011000011001100001100110000110011000011001100001100110000110;
        boldCharacters[78] = 200'b0110000110011100011001110001100111000110011110011001111001100111100110011011011001101101100110110110011011011001100111100110011110011001111001100111100110000110;
        boldCharacters[79] = 200'b0011111100011111111001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011001111111100011111100;
        boldCharacters[80] = 200'b0111111000011111110001100001100110000110011000011001100001100111111100011111100001100000000110000000011000000001100000000110000000011000000001100000000110000000;
        boldCharacters[81] = 200'b0001111000001111110001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011001101001100110010110011000111000111111000001111010;
        boldCharacters[82] = 200'b0111111000011111110001100001100110000110011000011001100001100111111100011111100001110000000111100000011111000001100110000110001100011000110001100001100110000110;
        boldCharacters[83] = 200'b0001111000001111110001100001100110000110011000000001100000000111000000001111100000011111000000000110000000011000000001100110000110011000011000111111000001111000;
        boldCharacters[84] = 200'b0111111110011111111000011110000001111000000111100000011110000001111000000111100000011110000001111000000111100000011110000001111000000111100000011110000001111000;
        boldCharacters[85] = 200'b0110000110011000011001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011001100001100110000110011000011000111111000001111000;
        boldCharacters[86] = 200'b0110000110011000011001100001100110000110011000011001100001100011001100001100110000110011000011001100001100110000011110000001111000000111100000011110000000110000;
        boldCharacters[87] = 200'b0110000110011000011001100001100110000110011000011001100001100110000110011000011001100001100110110110011111111001111111100111001110011100111001110011100110000110;
        boldCharacters[88] = 200'b0110000110011000011000110011000011001100000111100000011110000001111000000011000000001100000001111000000111100000011110000011001100001100110001100001100110000110;
        boldCharacters[89] = 200'b0110000110011000011000110011000011001100000111100000011110000001111000000011000000001100000000110000000011000000001100000000110000000011000000001100000000110000;
        boldCharacters[90] = 200'b0111111110011111111000000001100000001100000000110000000110000000011000000011000000001100000001100000000110000000110000000011000000011000000001111111100111111110;

        italicCharacters[65] = 200'b0000000110000000100100000110010000010001000010000100001000100000100010000100011000111111000010000100011000010001000001000100000100100000010010000010001000001000;
        italicCharacters[66] = 200'b0011111110001000000100100000010010000001001000000101100000010100000010010000001001111111000100000010010000001011000000101000000010100000010010000001001111111000;
        italicCharacters[67] = 200'b0000111111000100000000100000000010000000001000000001000000000100000000010000000001000000001000000000100000000010000000001000000000100000000001000000000011111100;
        italicCharacters[68] = 200'b0011111100001000001000100000010010000001001000000101000000010100000001010000001001000000100100000010100000001010000000101000000010100000010010000010001111110000;
        italicCharacters[69] = 200'b0001111111001000000000100000000010000000001000000001000000000100000000011111110001000000000100000000100000000010000000001000000000100000000010000000001111111000;
        italicCharacters[70] = 200'b0001111111001000000000100000000010000000001000000001000000000111111100010000000001000000000100000000100000000010000000001000000000100000000010000000001000000000;
        italicCharacters[71] = 200'b0000111111000100000000100000000010000000001000000000100000000100000000010000000001000011100100000010100000010010000001001000001000100000100010000010000111111000;
        italicCharacters[72] = 200'b0010000001001000000100100000010010000001001000000101000000100100000010011111111001000000100100000010100000010010000001001000000100100000010010000001001000000100;
        italicCharacters[73] = 200'b0011111111000001100000000110000000011000000001100000001100000000110000000011000000001100000000110000000110000000011000000001100000000110000000011000001111111100;
        italicCharacters[74] = 200'b0000111111000000000100000000010000000001000000000100000000010000000001000000001000000000100000000010000000010000000001000000000100100000010010000010000111110000;
        italicCharacters[75] = 200'b0010000010001000001000100000100100000100010000100001000010000100010000011110000001000100000100010000100000100010000010001000001000100000100010000010001000001000;
        italicCharacters[76] = 200'b0010000000001000000000100000000010000000001000000001000000000100000000010000000001000000000100000000100000000010000000001000000000100000000010000000001111111100;
        italicCharacters[77] = 200'b0011000011001010010100101001010010011001001001100101000000100100000010010000001001000000100100000010100000010010000001001000000100100000010010000001001000000100;
        italicCharacters[78] = 200'b0011000001001010000100101000010010100001001010000101000100100100010010010001001001000100100100010010100001010010000101001000010100100001010010000101001000001100;
        italicCharacters[79] = 200'b0001111110001000000100100000010010000001001000000101000000100100000010010000001001000000100100000010100000010010000001001000000100100000010010000001000111111000;
        italicCharacters[80] = 200'b0011111100001000001000100000010010000001001000000101000000100100000100011111100001000000000100000000100000000010000000001000000000100000000010000000001000000000;
        italicCharacters[81] = 200'b0000111100000100001000100000010010000001001000000101000000100100000010010000001001000000100100000010100010010010001001001000010100100001010001000010000011110100;
        italicCharacters[82] = 200'b0011111100001000001000100000010010000001001000000101000000100100000100011111100001000000001011000000100010000010000100001000010000100000100010000010001000001000;
        italicCharacters[83] = 200'b0000011100000110001000100000010010000001001000000000100000000010000000000111100000000001100000000010000000001000000001001000000100100000010001000010000011110000;
        italicCharacters[84] = 200'b0011111111000001100000000110000000011000000001100000001100000000110000000011000000001100000000110000000110000000011000000001100000000110000000011000000001100000;
        italicCharacters[85] = 200'b0010000001001000000100100000010010000001001000000101000000100100000010010000001001000000100100000010100000010010000001001000000100100000010001000010000011110000;
        italicCharacters[86] = 200'b0001000001000100000100010000010001000001000100000100100000100010000100001000010000100001000010000100001000100001000100000100010000010001000001001000000011000000;
        italicCharacters[87] = 200'b0010000001001000000100100000010010000001001000000101000000100100000010010000001001000000100100000010100110010010011001001010010100101001010010100101001100001100;
        italicCharacters[88] = 200'b0001000001000100000100001000100000100010000010010000010010000001001000000011000000001100000001001000001000100000100010000100001000010000010010000001001000000100;
        italicCharacters[89] = 200'b0010000001001000000100010000100001000010000100010000010010000001001000000011000000001100000000110000000110000000011000000001100000000110000000011000000001100000;
        italicCharacters[90] = 200'b0011111111000000000100000000100000000100000000010000000010000000010000000010000000001000000001000000001000000001000000000100000000100000000010000000001111111100;

        boldItalicCharacters[65] = 200'b0000000110000000111100000111110000011011000011001100001101100000110110000111111000111111000011001100011100110001100011000110001100110000110011000110001100011000;
        boldItalicCharacters[66] = 200'b0011111110001100001100110000110011000011001100001101110000110110000110011111111001111111000110000110011000011011100001101100000110110000010011000011001111111000;
        boldItalicCharacters[67] = 200'b0000111111000111111100110000000011000000001100000001100000000110000000011000000001100000001100000000110000000011000000001100000000110000000001111111000011111100;
        boldItalicCharacters[68] = 200'b0011111100001111111000110000110011000011001100001101100000110110000011011000011001100001100110000110110000011011000001101100000110110000110011111110001111110000;
        boldItalicCharacters[69] = 200'b0001111111001111111100110000000011000000001100000001100000000110000000011111110001111111000110000000110000000011000000001100000000110000000011111110001111111000;
        boldItalicCharacters[70] = 200'b0001111111001111111100110000000011000000001100000001100000000111111100011111110001100000000110000000110000000011000000001100000000110000000011000000001100000000;
        boldItalicCharacters[71] = 200'b0000111111000111111100110000000011000000001100000000110000000110000000011000111001100011100110000110110000110011000011001100011000110001100011111110000111111000;
        boldItalicCharacters[72] = 200'b0011000011001100001100110000110011000011001100001101100001100110000110011111111001111111100110000110110000110011000011001100001100110000110011000011001100001100;
        boldItalicCharacters[73] = 200'b0011111111001111111100001111000000111100000011110000011110000001111000000111100000011110000001111000001111000000111100000011110000001111000011111111001111111100;
        boldItalicCharacters[74] = 200'b0000111111000011111100000000110000000011000000001100000000110000000011000000011000000001100000000110000000110000000011000000001100110000110011111110000111110000;
        boldItalicCharacters[75] = 200'b0011000110001100011000110001100110001100011001100001100110000111110000011110000001101100000110110000110001100011000110001100011000110001100011000110001100011000;
        boldItalicCharacters[76] = 200'b0011000000001100000000110000000011000000001100000001100000000110000000011000000001100000000110000000110000000011000000001100000000110000000011111111001111111100;
        boldItalicCharacters[77] = 200'b0011000011001110011100111001110011111101001111110101100110110110000110011000011001100001100110000110110000110011000011001100001100110000110011000011001100001100;
        boldItalicCharacters[78] = 200'b0011000011001110001100111000110011100011001110001101101101100110110110011011011001101101100110110110110011110011001111001100111100110011110011001111001100011100;
        boldItalicCharacters[79] = 200'b0001111110001111111100110000110011000011001100001101100001100110000110011000011001100001100110000110110000110011000011001100001100110000110011111111000111111000;
        boldItalicCharacters[80] = 200'b0011111100001111111000110000110011000011001100001101100001100111111100011111100001100000000110000000110000000011000000001100000000110000000011000000001100000000;
        boldItalicCharacters[81] = 200'b0000111100000111111000110000110011000011001100001101100000100110000110011000011001100001100110000110110011011011001101001100011100110001100001111111000011101100;
        boldItalicCharacters[82] = 200'b0011111100001111111000110000110011000011001100001101110001100111111100011111100001100000001111000000111110000011001100001100110000110001100011000110001100011000;
        boldItalicCharacters[83] = 200'b0000011100000111111000111000110011000011001100000000110000000011000000000111100000011111100000000110000000011000000011001100001100110000110001111110000011110000;
        boldItalicCharacters[84] = 200'b0011111111001111111100001111000000111100000011110000011110000001111000000111100000011110000001111000001111000000111100000011110000001111000000111100000011110000;
        boldItalicCharacters[85] = 200'b0011000011001100001100110000110011000011001100001101100001100110000110011000011001100001100110000110110000110011000011001100001100110000110001111110000011110000;
        boldItalicCharacters[86] = 200'b0001100011000110001100011000110001100011000110001100110001100011001100001100110000110011000011001100001101100001101100000110110000011011000001111000000011000000;
        boldItalicCharacters[87] = 200'b0011000011001100001100110000110011000011001100001101100001100110000110011000011001100001100110000110110110110011011011001111111100111001110011100111001100001100;
        boldItalicCharacters[88] = 200'b0001100011000110001100001101100000110110000011010000011010000001101000000011000000001100000001111000001101100000110110000110011000011000110011000011001100001100;
        boldItalicCharacters[89] = 200'b0011000011001100001100011001100001100110000110110000011110000001111000000011000000001100000000110000000111000000011000000001100000000110000000011000000001100000;
        boldItalicCharacters[90] = 200'b0011111111001111111100000000110000000110000000011000000011000000011000000011000000001100000001100000001100000001100000000110000000110000000011111111001111111100;    end

    /*********************
     **     COUNTER     **
     *********************/
    reg [9:0] hCount = 0;
    reg [9:0] vCount = 0;

    wire hDisp = H_BPORCH <= hCount && hCount < H_BPORCH + H_VISIBLE;
    wire vDisp = V_BPORCH <= vCount && vCount < V_BPORCH + V_VISIBLE;
    wire hSync = H_BPORCH + H_VISIBLE + H_FPORCH <= hCount && hCount <= H_END;
    wire vSync = V_BPORCH + V_VISIBLE + V_FPORCH <= vCount && vCount <= V_END;

    reg [5:0] charX = 0;
    reg [4:0] charY = 0;
    reg [3:0] charU = 0;
    reg [4:0] charV = 0;

    always @(posedge VGA_CLK)
    begin
    	// NEW LINE
    	if (hCount == H_END)
    	begin
    		hCount <= 0;
    		charX <= 0;
    		charU <= 0;

    		// NEW FRAME
    		if (vCount == V_END)
    		begin
    			vCount <= 0;
    			charY <= 0;
    			charV <= 0;
    		end
    		// MID FRAME
    		else
    		begin
    			vCount <= vCount + 1;

                // end of BP; align charV and charY to 0
                if (vCount == V_BP_END) begin
                    charV <= 0;
                    charY <= 0;
                end
                else begin
                    // END CHAR
                    if (charV == 19)
                    begin
                        charV <= 0;
                        charY <= charY + 1;
                    end
                    // MID CHAR
                    else
                    begin
                        charV <= charV + 1;
                    end
                end
    		end
    	end
    	// MID LINE
    	else
    	begin
    		hCount <= hCount + 1;

            // end of BP; align charU and charX to 0
            if (hCount == H_BP_END) begin
                charU <= 0;
                charX <= 0;
            end
            else begin
                // END CHAR
                if (charU == 9)
                begin
                    charU <= 0;
                    charX <= charX + 1;
                end
                // MID CHAR
                else
                begin
                    charU <= charU + 1;
                end
            end
    	end
    end


    wire [10:0] wrAddr = charWrX | charWrY << 6;
    wire [10:0] readAddr = charX | charY << 6;
    wire [63:0] vramOut;
    RAM #(11, 64, 1) vram (
        .clk(CLOCK_50),

        .address_a(wrAddr),
        .wren_a(charWr),
        .data_a({charWrFlags, charWrFgColor, charWrBgColor, charWrCode}),
        .rden_a(1'b0),
        .q_a(),

        .address_b(readAddr),
        .wren_b(1'b0),
        .data_b(32'b0),
        .rden_b(1'b1),
        .q_b(vramOut)
    );

    wire [0:159] character = bold && italic
        ? boldItalicCharacters[vramOut[7:0]]
        : bold ? boldCharacters[vramOut[7:0]]
        : italic ? italicCharacters[vramOut[7:0]]
        : characters[vramOut[7:0]];
    wire [159:0] rvsCharacter = character;

    wire [0:9] line = charV < 16
        ? strikethrough && charV == 7 ? 10'h3FF : flipVertical ? rvsCharacter[charV*10 +: 10] : character[charV*10 +: 10]
        : underlined && charV == 17 ? 10'h3FF : 10'b0;
    wire [9:0] rvsLine = line;

    wire [23:0] color = (flipHorizontal ? rvsLine[charU] : line[charU]) ? vramOut[55:32] : vramOut[31:8];
    wire bold = vramOut[56];
    wire italic = vramOut[57];
    wire underlined = vramOut[58];
    wire strikethrough = vramOut[59];
    wire flipHorizontal = vramOut[60];
    wire flipVertical = vramOut[61];

    assign VGA_HS = ~hSync;
    assign VGA_VS = ~vSync;
    assign VGA_R = ~VGA_BLANK_N ? 0 : color[23:16];
    assign VGA_G = ~VGA_BLANK_N ? 0 : color[15:8];
    assign VGA_B = ~VGA_BLANK_N ? 0 : color[7:0];
    assign VGA_BLANK_N = ~(~hDisp || ~vDisp);
    assign VGA_SYNC_N = ~(hSync ^ vSync);
endmodule